/* This version uses num_real_pages and num_real_patterns */
/*
 * pattern: 12-bit
 * (12-bit)comparator*32ea for one block (384-bit)
 * Total 128 blocks array (384*128=49152-bit)
 *
 * 4096 * 12 = 49152
 * PPB=64, NOB=64, NOP=4096
 */

`define NOP 4096 // total number of pages // 4096
`define P_SIZE 12 // number of bits in pattern (=number of bits in page)
`define ARR_SIZE ((`NOP)*(`P_SIZE)) // number of bits in input array (4096 page * 12-bit) // 49152

`define PPB 64 // number of page comparators per block
`define NOB ((`NOP)/(`PPB)) // number of blocks (=comparing epoch) // 64
//`define B_SIZE (`ARR_SIZE)/(`NOB) // number of bits in a block // 768
`define B_SIZE 768 // Velog must determine specific number of bits for assignment

`define NOP_WIDTH 12 // integer which can store the range of page number 0~4095 (12-bit can store 0~4095 integer)
`define NOB_WIDTH 6 // integer which can store the range of block number 0~63 (6-bit can store 0~63 integer)
`define PPB_WIDTH 6 // integer which can store the range of block number 0~63 (6-bit can store 0~63 integer)

`define B_OFS_WIDTH 10 // integer which can store the range of block offset(in-block bit index) 0~768(=0 ~ NOP_WIDTH*PPB) (10-bit can store 0~1023)

`define MAX_TPN_NUM 8 // number of true pages are from 1 to 8
`define MAX_TPN_NUM_WIDTH 4 // integer which can store the range of max tpn number 0~8 (4-bit can store 0~15)

`define NUM_PATT_WIDTH 3 // integer which can store 000, 001, 011, 111 and 1~4 (3-bit can store 0~7)

/*
 * One comparator can compare one page with four page-size patterns
 * In one epoch, HW finds true pages which are equal to patterns in one block
 * After processing all blocks, HW returns an array which consists of the index number of true pages
 */

/* testbench.sv */

module find_bit_pattern_tb;
  // Inputs
  reg clk;
  reg rst;
  reg [`B_SIZE-1:0] arr;
  reg [`P_SIZE-1:0] pattern1, pattern2, pattern3, pattern4;
  reg [`NOB_WIDTH:0] block_index;
  reg put_global;
  
  // New inputs
  integer num_real_pages;
  reg [2:0] num_real_patterns;
  
  integer num_real_blocks;
   
  // Outputs
  reg [`MAX_TPN_NUM*`NOP_WIDTH-1:0] tpn_arr;
  reg [`MAX_TPN_NUM_WIDTH-1:0] num_truepages;
  
  integer i;
  
  top f1
  (
    .out(tpn_arr),
    .num_tpn(num_truepages),
    .clk(clk),
    .rst(rst),
    .b_idx(block_index),
    .a(arr),
    .x1(pattern1),
    .x2(pattern2),
    .x3(pattern3),
    .x4(pattern4),
    .put_global_array(put_global),
    .num_real_patterns(num_real_patterns)
  );
  
  initial begin
    forever
      #10 clk = ~clk;
  end
  
  initial begin
    #50
    forever begin
      put_global = 1;
      #10
      put_global = 0;
      #30
      put_global = 0;
    end
  end
  
  //`define BASIC
  initial
    begin
      $dumpfile("top.vcd");
      $dumpvars(2,f1);
      // Initialize Inputs
      clk = 1'b0;
      rst = 1'b0;
      put_global = 0;
      #10 
      
      rst = 1'b1;
      pattern2 = 12'h111;
      pattern1 = 12'h232;
      pattern3 = 12'h333;
      pattern4 = 12'h444;
      
      // Start
      block_index = `NOB_WIDTH'd0;
      
      /* Maximum 4096 pages(12-bit binary-encoded) (called page in this verilog code) */
      `ifdef BASIC
        $display("number of real page is set to 4096");
        num_real_pages = `NOP_WIDTH'd4095;
      	num_real_patterns = 3'd4;
      `endif
      `ifndef BASIC
        $display("number of real page is different with 4096");
        num_real_pages = `NOP_WIDTH'd4095;
      	num_real_patterns = 3'd3;
      `endif
      
      num_real_blocks = num_real_pages / `NOB;
      for (i=1; i<=num_real_blocks; i=i+1) begin
        #40
        block_index = block_index+1;
      end
      #40
      block_index = block_index+1;
      
      #40
      rst = 1'b0;
      
      #20 $finish;
      
    end
  
  /* input vector array with block unit */
  // Expected output: 2, 40, 5e, 7e, 140, 145, 165, fc2
  initial begin
    #10
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_111_222_222;
    #40
    arr = `B_SIZE'h222_333_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_333_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_333;
    #40
    arr = `B_SIZE'h666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_999;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_888;
    #40
    
    arr = `B_SIZE'h555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_222_222_111_555_555_555_555_555__555_555_555_222_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_555_222_222_111_555_555_555_555_333;
    #40
    
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_444;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_555;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_444_666;
    #40
    arr = `B_SIZE'h222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_222_333_222_555;
    //#40
  end
 
endmodule // find_bit_pattern_tb
